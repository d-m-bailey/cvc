.INCLUDE lib.cdl
.INCLUDE "lib.cdl"
.INCLUDE $CDL_PATH/lib.cdl
.INCLUDE "$CDL_PATH/lib.cdl"


.SUBCKT TOP P1 P2
X1 P1 P2 res
X2 P1 P2 res2
.ENDS


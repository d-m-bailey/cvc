.SUBCKT res POS NEG
R0 POS NET 10.0
.ENDS
.SUBCKT res2 POS NEG
R0 POS NET 20.0
.ENDS
